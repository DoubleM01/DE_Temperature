`timescale 1ns/1ps 
module temp_tb ();  
reg clk, rst; 
wire 