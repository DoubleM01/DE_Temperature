module lcd(
    clk,
    e
);