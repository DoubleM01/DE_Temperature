module lcd();